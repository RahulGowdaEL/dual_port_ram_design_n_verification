package mem_package;
    import uvm_pkg::*;
   `include "uvm_macros.svh"
   `include "mem_seqr.sv"
   `include "mem_driver.sv"
   `include "mem_monitor.sv"
   `include "mem_seq_item.sv"
   `include "mem_sequence.sv"
   `include "mem_agent.sv"
   `include "mem_wr_rd_test.sv"
   `include "mem_env.sv"
   `include "mem_soreboard"
   `include "tb_top.sv"
endpackage
